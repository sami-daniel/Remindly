module main

import database

type UnitOfWork = database.UnitOfWork

fn main() {
	
}